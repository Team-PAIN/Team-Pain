`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:50:49 11/27/2012 
// Design Name: 
// Module Name:    localization 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module localization(
		output [7:0] ANGLE,
		output [1:0] ANGLE_DIRECTION,
		output [7:0] DISTANCE1,
		output [7:0] DISTANCE2
    );


endmodule
